library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY prac8 IS

PORT	(CLK, BOTON, RX: IN STD_LOGIC;
		TX:		OUT STD_LOGIC;
		SWITCH:	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DOUT:		OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END prac8;

ARCHITECTURE Behavioral OF prac8 IS

COMPONENT RS232 IS
GENERIC	(FPGA_CLK:		INTEGER;
			BAUD_RS232:	INTEGER);
PORT		(CLK:		IN STD_LOGIC;
			RX:		IN STD_LOGIC;
			TX_INI:	IN STD_LOGIC;
			TX_FIN:	OUT STD_LOGIC;
			TX:		OUT STD_LOGIC;
			RX_IN:	OUT STD_LOGIC;
			DATAIN:	IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			DOUT:		OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

SIGNAL TX_INI_S, TX_FIN_S, RX_IN_S: STD_LOGIC;
SIGNAL DATAIN_S, DOUT_S, midato: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL SWITCHTEST: STD_LOGIC_VECTOR(3 DOWNTO 0):="0011";

BEGIN

recepcion: PROCESS(CLK, RX_IN_S)
BEGIN
	IF RISING_EDGE(CLK) THEN
		IF (RX_IN_S='1') THEN
			DOUT <= std_logic_vector(unsigned(DOUT_S(7 DOWNTO 0))-48)(3 downto 0);
		END IF;
	END IF;
END PROCESS;

transmision: PROCESS(CLK)
BEGIN
	IF RISING_EDGE(CLK) THEN
		DATAIN_S <= std_logic_vector(unsigned(("0000"& SWITCH))+48);
	END IF;
END PROCESS;

TX_INI_S <= NOT BOTON;

UART: RS232
GENERIC MAP(
	FPGA_CLK => 12000000,	--FRECUENCIA DEL FPGA 
	BAUD_RS232 => 9600		--BAUDIOS
)
PORT MAP(
	CLK => CLK,
	RX => RX,
	TX_INI => TX_INI_S,
	TX_FIN => TX_FIN_S,
	TX => TX,
	RX_IN => RX_IN_S,
	DATAIN => DATAIN_S,
	DOUT => DOUT_S
);

END Behavioral;